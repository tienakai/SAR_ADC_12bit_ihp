** sch_path: /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.tech/xschem/sg13g2_tests_xyce/dc_hv_pmos.sch
**.subckt dc_hv_pmos
Vgs GND net1 0
Vds GND net3 0
XM1 GND net1 net2 GND sg13_hv_pmos w=1.0u l=0.45u ng=1 m=1
Vd net2 net3 0
.save i(vd)
**** begin user architecture code







.lib cornerMOShv.lib mos_tt





.param temp=27
.control
save all
dc Vds 0 3.0 0.01 Vgs 0.3 1.5 0.05
write dc_hv_pmos.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
