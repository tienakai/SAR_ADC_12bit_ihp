** sch_path: /home/tien/ihp/schematic/simulations/bootstrap_tb.sch
**.subckt bootstrap_tb
x1 VDD VGATE VSS SW_ON VIN EN bootstrap
V9 EN VSS pulse(0 1.8 0 0.1n 0.1n 50n 100n)
V13 VIN VSS sin(0.6 0.6 100k 0 0 0)
V1 VDD VSS 1.8
.save i(v1)
V4 VSS GND 0
C1 VIN_SMPL VSS 2p m=1
XM1 VIN_SMPL VGATE VIN VSS sg13_lv_nmos w=17u l=0.13u ng=4 m=1
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.include /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice




.option temp = 27
.save all

.option GMIN=1e-12 reltol=1e-6

.tran 10n 100u


**** end user architecture code
**.ends

* expanding   symbol:  bootstrap/bootstrap.sym # of pins=6
** sym_path: /home/tien/ihp/schematic/bootstrap/bootstrap.sym
** sch_path: /home/tien/ihp/schematic/bootstrap/bootstrap.sch
.subckt bootstrap VDD VGATE VSS SW_ON VIN EN
*.ipin VDD
*.ipin VSS
*.ipin VIN
*.ipin EN
*.opin VGATE
*.opin SW_ON
XM5 VDD VGATE Vtop Vtop sg13_lv_pmos w=0.32u l=0.15u ng=1 m=1
XM1 VGATE EN_Z_LVL_SHFT Vtop Vtop sg13_lv_pmos w=16u l=0.38u ng=4 m=1
XM2 Vtop Vbottom Vtop Vtop sg13_lv_pmos w=10u l=10u ng=2 m=1
XM6 EN_Z_LVL_SHFT EN VDD VDD sg13_lv_pmos w=0.35u l=0.15u ng=1 m=1
XM7 EN_Z_LVL_SHFT EN Vbottom VSS sg13_lv_nmos w=0.63u l=0.15u ng=1 m=1
XM8 EN_Z_LVL_SHFT VGATE Vbottom VSS sg13_lv_nmos w=1.8u l=0.15u ng=2 m=1
XM3 Vbottom EN_Z VSS VSS sg13_lv_nmos w=3.5u l=0.15u ng=1 m=1
XM10 VIN VGATE Vbottom VSS sg13_lv_nmos w=3.5u l=0.15u ng=1 m=1
XM4 net2 EN_Z VSS VSS sg13_lv_nmos w=3.5u l=0.15u ng=1 m=1
XM11 VGATE VDD VGATE_1V8 VSS sg13_lv_nmos w=3.5u l=0.45u ng=1 m=1
XM9 VGATE VDD net2 VSS sg13_hv_nmos w=6.3u l=0.45u ng=2 m=1
x2 SW_ON net1 VDD VSS sg13g2_inv_2
x4 net1 VGATE_1V8 VDD VSS sg13g2_inv_1
x1 EN_Z EN VDD VSS sg13g2_inv_1
.ends

.end
