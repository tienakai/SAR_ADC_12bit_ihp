** sch_path: /home/tien/ihp/schematic/simulations/latch_comparator_tb2.sch
**.subckt latch_comparator_tb2
x1 VDD vinp Vbias outp clk outm GND latched_comparator
V1 VDD GND 1.2
V5 Vbias GND DC 1
V6 clk GND PULSE(0 1.2 0 1n 1n 5n 100n)
V8 vinp GND DC 1.05
C1 Vbias GND 6.4p m=1
C4 outp GND 50f m=1
C2 vinp GND 6.4p m=1
C3 outm GND 50f m=1
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.include /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27
.param clock = 100e6       ; 100 MHz clock
.param period = {1/clock}
.param num_cycles = 100
.param tr = {num_cycles * period}

.control
save all
* Operating point simulation
op

set appendwrite

* Transient analysis
.options meas_step_max=1e-10
tran 500p 1u
let vindiff = v(vinp) - v(vbias)
let clk = v(clk)
let vout = v(outp) - v(outm)

meas TRAN rise_time TRIG v(outp) VAL=0.12  TD=9n RISE=4 TARG v(outp) VAL=1.08 TD=9n RISE=4
meas TRAN fall_time TRIG v(outp) VAL=1.08  TD=9n RISE=4 TARG v(outp) VAL=0.12 TD=9n RISE=4


.endc


**** end user architecture code
**.ends

* expanding   symbol:  latched_comparator/latched_comparator.sym # of pins=7
** sym_path: /home/tien/ihp/schematic/latched_comparator/latched_comparator.sym
** sch_path: /home/tien/ihp/schematic/latched_comparator/latched_comparator.sch
.subckt latched_comparator VDD Vin_P Vin_N OUT_P EN OUT_N VSS
*.ipin Vin_P
*.ipin Vin_N
*.iopin VDD
*.iopin VSS
*.ipin EN
*.opin OUT_P
*.opin OUT_N
XM1 net1 ENi VDD VDD sg13_lv_pmos w=0.32u l=0.15u ng=1 m=1
XM2 OUT_Ni ENi VDD VDD sg13_lv_pmos w=0.32u l=0.15u ng=1 m=1
XM3 OUT_Ni OUT_Pi VDD VDD sg13_lv_pmos w=1.25u l=0.15u ng=1 m=1
XM4 net2 ENi VDD VDD sg13_lv_pmos w=0.32u l=0.15u ng=1 m=1
XM5 OUT_Pi ENi VDD VDD sg13_lv_pmos w=0.32u l=0.15u ng=1 m=1
XM6 OUT_Pi OUT_Ni VDD VDD sg13_lv_pmos w=1.25u l=0.15u ng=1 m=1
XM7 net1 Vin_P net3 VSS sg13_lv_nmos w=0.55u l=0.13u ng=1 m=1
XM8 net2 Vin_N net3 VSS sg13_lv_nmos w=0.55u l=0.13u ng=1 m=1
XM9 OUT_Pi OUT_Ni net2 VSS sg13_lv_nmos w=0.42u l=0.15u ng=1 m=1
XM10 OUT_Ni OUT_Pi net1 VSS sg13_lv_nmos w=0.42u l=0.15u ng=1 m=1
XM11 net3 net3 net3 VSS sg13_lv_nmos w=0.55u l=0.13u ng=1 m=2
XM12 net3 ENi VSS VSS sg13_lv_nmos w=0.9u l=0.15u ng=1 m=2
x4 net4 OUT_Pi VDD VSS sg13g2_inv_2
x5 net5 OUT_Ni VDD VSS sg13g2_inv_2
x1 ENi EN VDD VSS sg13g2_buf_4
x6 OUT_P net4 VDD VSS sg13g2_inv_4
x2 OUT_N net5 VDD VSS sg13g2_inv_4
.ends

.GLOBAL VDD
.GLOBAL GND
.end
