** sch_path: /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/iso_dc_lv_nmos.sch
**.subckt iso_dc_lv_nmos
Vgs G S 1.2
Vds D S 1.5
Vd D net1 0
.save i(vd)
XM1 net1 G S iso_B sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XD1 S net2 sub! isolbox l=10.0u w=10.0u
XR1 GND sub! ptap1 R=262.8 w=0.78e-6 l=0.78e-6
XR2 S iso_B ptap1 R=262.8 w=0.78e-6 l=0.78e-6
Vdd net2 GND 1.5
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.include diodes.lib



.param temp=27
.control
save all
op
write iso_dc_lv_nmos.raw
set appendwrite
dc Vds 0 1.2 0.01 Vgs 0.3 1.0 0.1
write iso_dc_lv_nmos.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL sub!
.end
