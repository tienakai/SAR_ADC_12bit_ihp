** sch_path: /home/tien/ihp/schematic/simulations/latched_comparator_tb.sch
**.subckt latched_comparator_tb
x1 VDD inp inn OUT_P EN_COMP OUT_N GND latched_comparator
V1 VDD GND 1.8
V3 inp GND 0 PULSE(1.2 1.3 0 0.1n 0.1n 80n 200n)
V2 inn GND 0 PULSE(1.3 1.2 0 0.1n 0.1n 80n 200n)
V7 EN_COMP GND 0 PULSE(0 1.8 0 0.1n 0.1n 50n 100n)
.save i(v7)
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.include /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice




.option temp = 27
.save all

.option GMIN=1e-12 reltol=1e-6

.tran 10n 100u


**** end user architecture code
**.ends

* expanding   symbol:  latched_comparator/latched_comparator.sym # of pins=7
** sym_path: /home/tien/ihp/schematic/latched_comparator/latched_comparator.sym
** sch_path: /home/tien/ihp/schematic/latched_comparator/latched_comparator.sch
.subckt latched_comparator VDD Vin_P Vin_N OUT_P EN OUT_N VSS
*.ipin Vin_P
*.ipin Vin_N
*.iopin VDD
*.iopin VSS
*.ipin EN
*.opin OUT_P
*.opin OUT_N
XM1 net1 ENi VDD VDD sg13_lv_pmos w=0.32u l=0.15u ng=1 m=1
XM2 OUT_Ni ENi VDD VDD sg13_lv_pmos w=0.32u l=0.15u ng=1 m=1
XM3 OUT_Ni OUT_Pi VDD VDD sg13_lv_pmos w=1.25u l=0.15u ng=1 m=1
XM4 net2 ENi VDD VDD sg13_lv_pmos w=0.32u l=0.15u ng=1 m=1
XM5 OUT_Pi ENi VDD VDD sg13_lv_pmos w=0.32u l=0.15u ng=1 m=1
XM6 OUT_Pi OUT_Ni VDD VDD sg13_lv_pmos w=1.25u l=0.15u ng=1 m=1
XM7 net1 Vin_P net3 VSS sg13_lv_nmos w=0.55u l=0.13u ng=1 m=1
XM8 net2 Vin_N net3 VSS sg13_lv_nmos w=0.55u l=0.13u ng=1 m=1
XM9 OUT_Pi OUT_Ni net2 VSS sg13_lv_nmos w=0.42u l=0.15u ng=1 m=1
XM10 OUT_Ni OUT_Pi net1 VSS sg13_lv_nmos w=0.42u l=0.15u ng=1 m=1
XM11 net3 net3 net3 VSS sg13_lv_nmos w=0.55u l=0.13u ng=1 m=2
XM12 net3 ENi VSS VSS sg13_lv_nmos w=0.9u l=0.15u ng=1 m=2
x4 net4 OUT_Pi VDD VSS sg13g2_inv_2
x5 net5 OUT_Ni VDD VSS sg13g2_inv_2
x1 ENi EN VDD VSS sg13g2_buf_4
x6 OUT_P net4 VDD VSS sg13g2_inv_4
x2 OUT_N net5 VDD VSS sg13g2_inv_4
.ends

.GLOBAL GND
.GLOBAL VDD
.end
