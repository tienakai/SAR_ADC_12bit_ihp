** sch_path: /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/inv_mc_tb.sch
**.subckt inv_mc_tb
VDD1 vdd GND 1.5
XM1 inv_out inv_in GND GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 inv_out inv_in vdd vdd sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM3 GND inv_out GND GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
VIN1 in GND dc 0.75 ac 1 sin(0.75 1m 100Meg)
R1 inv_out inv_in 100Meg m=1
XC1 inv_in in cap_cmim w=10.0e-6 l=10.0e-6 m=7
**** begin user architecture code


** IHP models
.lib cornerMOSlv.lib mos_tt_stat
.lib cornerMOShv.lib mos_tt_stat
.lib cornerHBT.lib hbt_typ_stat
.lib cornerRES.lib res_typ_stat
.lib cornerCAP.lib cap_typ_stat





.control
set num_threads 1

ac dec 1001 1 100G
let gain_lin = abs(inv_out)
let gain_dB = vdb(inv_out)
meas ac gain_passband_dB max gain_dB
let gain_fc_dB = gain_passband_dB-3
meas ac fc_l when gain_dB = gain_fc_dB
meas ac fc_u when gain_dB = gain_fc_dB cross=last
let GBW = gain_lin[0] * (fc_u-fc_l)

echo results_save_begin
print gain_passband_dB
print fc_l
print fc_u
print GBW
echo results_save_end

.endc




**nr_workers=50
**nr_mc_sims=1000

**results_plot_begin
**gain_passband_dB
**fc_l
**fc_u
**GBW
**results_plot_end


**** end user architecture code
**.ends
.GLOBAL GND
.end
