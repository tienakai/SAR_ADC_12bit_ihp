** sch_path: /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.tech/xschem/sg13g2_tests_xyce/dc_lv_nmos.sch
**.subckt dc_lv_nmos
Vgs net1 GND 0.0
Vds net3 GND 0
Vd net3 net2 0
XM2 net2 net1 GND GND sg13_lv_nmos w=1.0u l=0.13u ng=1
**** begin user architecture code



.preprocess replaceground true
.option temp=27
.step  vgs 0.0 0.8 0.05
.dc vds 0 1.2 0.01
.print dc format=raw file=dc_lv_nmos.raw i(Vd)





.lib /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.tech/xyce/models/cornerMOSlv.lib mos_tt






**** end user architecture code
**.ends
.GLOBAL GND
.end
