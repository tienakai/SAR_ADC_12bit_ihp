** sch_path: /home/tien/ihp/schematic/test3.sch
**.subckt test3
Vgs G GND 1.2
Vds D GND 1.8
Vd D net1 0
.save i(vd)
XM5 net1 G GND GND sg13_lv_nmos w=34u l=0.13u ng=4 m=1
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt




.param temp=27
.control
save all
op
write test3.raw
set appendwrite
dc Vds 0 1.8 0.01
write test3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
