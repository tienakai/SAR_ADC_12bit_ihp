** sch_path: /home/tien/ihp/schematic/individual_switches/switch_C8.sch
**.subckt switch_C8 VIN EN_VIN VREF_GND EN_VSS Cbtm VSS VREF EN_VREF_Z EN_VCM VCM VDD
*.ipin VIN
*.ipin EN_VIN
*.ipin VREF_GND
*.ipin EN_VSS
*.opin Cbtm
*.iopin VSS
*.ipin VREF
*.ipin EN_VREF_Z
*.ipin EN_VCM
*.ipin VCM
*.iopin VDD
XM1 VREF_GND EN_VSS Cbtm VSS sg13_lv_nmos w=3.45u l=0.13u ng=1 m=1
XM2 Cbtm EN_VREF_Z VREF VDD sg13_lv_pmos w=16u l=0.35u ng=2 m=1
XM3 VCM EN_VCM Cbtm VSS sg13_lv_nmos w=4.5u l=0.13u ng=1 m=1
XM5 VIN EN_VIN Cbtm VSS sg13_lv_nmos w=0.9u l=0.13u ng=1 m=1
**.ends
.end
