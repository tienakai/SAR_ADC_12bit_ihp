** sch_path: /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/dc_lv_nmos.sch
**.subckt dc_lv_nmos
Vgs G GND 1.2
Vds D GND 1.5
Vd D net1 0
.save i(vd)
XM1 net1 G GND GND sg13_lv_nmos w=1.0u l=0.45u ng=1 m=1
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt




.param temp=27
.control
save all
op
write dc_lv_nmos.raw
set appendwrite
dc Vds 0 1.2 0.01 Vgs 0.3 1.0 0.1
write dc_lv_nmos.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
