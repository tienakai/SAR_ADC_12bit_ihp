** sch_path: /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.tech/xschem/sg13g2_tests_xyce/ac_rfmim_cap.sch
**.subckt ac_rfmim_cap
V1 in GND dc 0 ac 1
R2 out GND 100k m=1
XC1 in out GND cap_rfcmim w=10.0e-6 l=10.0e-6 wfeed=5.0e-6
**** begin user architecture code







.lib cornerCAP.lib cap_typ
.lib cornerRES.lib res_typ





.param temp=27
.control
ac dec 1000 1e6 1e9
let mag=abs(out)
meas ac freq_at when mag = 0.707
let C = 1/(2*PI*freq_at*1e+5)
print C
write ac_mim_cap.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
