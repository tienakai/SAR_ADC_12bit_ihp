** sch_path: /home/tien/conda-gf180mcu-env/share/pdk/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/dc_ntap1.sch
**.subckt dc_ntap1
Vres Vcc net1 1.5
Vr Vcc net2 0
.save i(vr)
Vres2 GND net1 0
XR4 net2 net1 ntap1 R=225.8 w=1.0e-6 l=0.78e-6
XR5 net2 net1 ntap1 R=30.62 w=10.0e-6 l=1.0e-6
**** begin user architecture code



.lib cornerRES.lib res_typ





.param temp=27
.control
save all
op
print Vcc/I(Vr)
reset
dc Vres 0 3 0.01
write dc_ntap1.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
