** sch_path: /home/tien/ihp/schematic/test4.sch
**.subckt test4
Vgs net1 GND -1.2
Vds net3 GND -1.8
Vd net3 net2 0
.save i(vd)
XM1 GND net1 net2 GND sg13_lv_pmos w=128u l=0.35u ng=16 m=1
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt



.options savecurrents
.param temp=27
.control
save all
op
write test4.raw
set appendwrite
dc Vds 0 -1.8 -0.01
write test4.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
